module test;
  initial begin
    $display("Hello, Verilog World!");
    $finish;
  end
endmodule